module AND(input wire a, input wire b, input wire c, output wire sum);
assign sum = a & b & c;
endmodule
